`ifndef FUNCTIONS_VH
`define FUNCTIONS_VH

function integer max(input integer a, input integer b);
    max = (a > b) ? a : b;
endfunction

`endif